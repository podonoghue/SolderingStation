*FDS4675 at Temp. Electrical Model
*----------------------------------
.SUBCKT FDS4675 20 10 30 50
*20=DRAIN 10=GATE 30=SOURCE 50=VTEMP
Rg 10 11x 1
Rdu 12x 1 1u
M1 2 1 4x 4x DMOS L=1u W=1u
.MODEL DMOS PMOS(VTO=-1.5 KP=6.33E+1
+THETA=.1 VMAX=9.5E5 LEVEL=3)
Cgs 1 5x 4220p
Rd 20 4 2.4E-3 
Dds 4 5x DDS
.MODEL DDS D(M=2.59E-1 VJ=2.48E-2 CJO=1568p)
Dbody 20 5x DBODY
.MODEL DBODY D(IS=1.75E-11 N=1.064513 RS=.00016 TT=16.08n)
Ra 4 2 2.4E-3 
Rs 5x 5 0.5m
Ls 5 30 0.5n
M2 1 8 6 6 INTER
E2 8 6 4 1 2
.MODEL INTER PMOS(VTO=0 KP=10 LEVEL=1)
Cgdmax 7 4 3450p
Rcgd 7 4 10meg
Dgd 4 6 DGD
Rdgd 4 6 10meg
.MODEL DGD D(M=1.58E-1 VJ=1.4E-6 CJO=3450p)
M3 7 9 1 1 INTER
E3 9 1 4 1 -2
*ZX SECTION
EOUT 4x 6x poly(2) (1x,0) (3x,0) 0 0 0 0 1
FCOPY 0 3x VSENSE 1
RIN 1x 0 1G
VSENSE 6x 5x 0
RREF 3x 0 10m
*TEMP SECTION
ED 101 0 VALUE {V(50,100)}
VAMB 100 0 25
EKP 1x 0 101 0 .005
*VTO TEMP SECTION
EVTO 102 0 101 0 .0015
EVT 11x 12x 102 0 1
*DIODE THEMO BREAKDOWN SECTION
EBL VB1 VB2 101 0 .08
VBLK VB2 0 40
D DB1 20 DBLK
.MODEL DBLK D(IS=1E-14 CJO=.1p RS=.1)
EDB 0 DB1 VB1 0 1
.ENDS FDS4675
*FDS4675 (Rev.B) 7/29/03 **ST

